library verilog;
use verilog.vl_types.all;
entity MaxAndar3_vlg_vec_tst is
end MaxAndar3_vlg_vec_tst;
