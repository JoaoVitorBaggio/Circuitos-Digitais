library verilog;
use verilog.vl_types.all;
entity INC8_vlg_vec_tst is
end INC8_vlg_vec_tst;
