library verilog;
use verilog.vl_types.all;
entity TopLevel_vlg_vec_tst is
end TopLevel_vlg_vec_tst;
