library verilog;
use verilog.vl_types.all;
entity Temporizador_vlg_vec_tst is
end Temporizador_vlg_vec_tst;
