library verilog;
use verilog.vl_types.all;
entity DEMUX1x8_vlg_vec_tst is
end DEMUX1x8_vlg_vec_tst;
