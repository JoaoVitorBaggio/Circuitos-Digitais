library verilog;
use verilog.vl_types.all;
entity FSM1_vlg_vec_tst is
end FSM1_vlg_vec_tst;
