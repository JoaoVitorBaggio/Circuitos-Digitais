library verilog;
use verilog.vl_types.all;
entity Compare3_vlg_vec_tst is
end Compare3_vlg_vec_tst;
