library verilog;
use verilog.vl_types.all;
entity Elevador_TL_vlg_vec_tst is
end Elevador_TL_vlg_vec_tst;
